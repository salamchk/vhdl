-------------------------------------------------------------------------------
--
-- Title       : 
-- Design      : lab2
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- File        : c:\My_Designs\lab2\compile\OR.vhd
-- Generated   : Sun Dec 13 00:12:45 2020
-- From        : c:\My_Designs\lab2\src\OR.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;

entity \OR\ is
  port(
       A : in STD_LOGIC_VECTOR(0 to 1);
       B : in STD_LOGIC_VECTOR(0 to 1);
       C : out STD_LOGIC_VECTOR(0 to 1)
  );
end \OR\;

architecture \OR\ of \OR\ is

begin

end \OR\;
